`timescale 1ps/1ps

module KECCAK_f_tb;

    // Inputs and Outputs
    logic [1599:0] S_in, S_out;
    
    // Instantiate the module under test
    KECCAK_p dut (
        .S_in(S_in),
        .S_out(S_out)
    );
    
    // Test stimulus
    initial begin
        // Apply stimulus
        S_in = 'h1F00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000008000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        //S_in = 'h000000000000001f_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_8000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000;
        
        // Wait for a few clock cycles
        #10;
        
        // Print the output
        $display("S_out =   %h", S_out);
        $display("Expected: 1E000000000000001F00000000000000000000000000008000000000000000003E0000000000000001000000000000001F00000000000000000000000000008000000000000000003E0000000000000001000000000000001F00000000000000000000000000008000000000000000003E0000000000000001000000000000001F00000000000080000000000000008000000000000000003E0000000000000001000000000000001F00000000000000000000000000008000000000000000003E00000000000000");
        
        // End the simulation
        $finish;
    end
    
endmodule
module pad (
    input [1087:0] data_in,
    input [10:0] data_length,
    output [1087:0] data_out,
    output [1087:0] data_next
);

    always_comb begin
        if ((data_length >= 0) && (data_length <= 1088)) begin
            if (data_length == 1088) begin
                data_out = data_in;
                data_next = 1088'b1f00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000008000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            end else if (data_length == 1087) begin
                data_out = {data_in[1088:8], 1'h1, data_in[7:1]};
                data_next = 1088'b0f00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000008000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            end else if (data_length == 1086) begin
                data_out = {data_in[1088:8], 2'h3, data_in[7:2]};
                data_next = 1088'b0700000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000008000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            end else if (data_length == 1085) begin
                data_out = {data_in[1088:8], 3'h7, data_in[7:3]};
                data_next = 1088'b0300000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000008000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            end else if (data_length == 1084) begin
                data_out = {data_in[1088:8], 4'hf, data_in[7:4]};
                data_next = 1088'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000008000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            end else if (data_length == 1083) begin
                data_out = {data_in[1088:8], 5'h1f, data_in[7:5]};
                data_next = 1088'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000008000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            end else if (data_length == 1082) begin
                data_out = {data_in[1088:8], 6'h3f, data_in[7:6]};
                data_next = 1088'b0;
            end else if (data_length == 1081) begin
                data_out = {data_in[1088:8], 7'b101_1111, data_in[7]};
                data_next = 1088'b0;
            end else if (data_length == 1080) begin
                data_out = {data_in[1088:8], 8'b1001_1111};
                data_next = 1088'b0;
            end else begin
                case (data_length % 8)
                    0: data_out = ;
                    1: data_out = ;
                    2: data_out = ;
                    3: data_out = ;
                    4: data_out = ;
                    5: data_out = ;
                    6: data_out = ;
                    7: data_out = ;
                    default: 
                endcase
                data_next = 1088'b0;
            end
        end else begin
            data_out = data_in;
            data_next = 1088'b0;            
        end
    end

endmodule
`timescale 1ps/1ps

module KECCAK_f_tb;

    logic [1599:0] S_in, S_out;
    logic clock, reset, done;
    
    KECCAK_f dut (.clock(clock), .reset(reset), .S_in(S_in), .S_out(S_out), .done(done));

    initial begin
        $dumpfile("KECCAK_f.vcd");
        $dumpvars;

        clock = 0;
        reset = 0;
      //S_in = 'h1F00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000008000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      //S_in = 'hF303000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000008000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      //S_in = 'ha3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a300000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        S_in = 'h53587bd907000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000008000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

        $display("S_in  = %h", S_in);
        $display;

        #1; reset = 1;
    end

    initial forever #1 clock = ~clock;

    initial begin
        repeat (24) begin
            #2;
            $display("Round %0d", $time/2);
            $display("S_out = %h", S_out);
            $display("Done  = %b", done);
            $display;
        end

	/*#1;
	S_in = S_out ^ 'h1f00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000008000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        $display("S_in  = %h", S_in);
        $display;

        repeat (25) begin
            #2;
            $display("Round %0d", $time/2);
            $display("S_out = %h", S_out);
            $display("Done  = %b", done);
            $display;
        end*/

	#1;
        $finish;
    end
    
endmodule

`timescale 1ps/1ps

module KECCAK_f_tb;

    // Inputs and Outputs
    //logic [1599:0] S_in, S_out;
    logic [63:0] A_in [0:4][0:4];
    logic [63:0] A_out [0:4][0:4];
    
    // Instantiate the module under test
    // KECCAK_f dut (
    //     .S_in(S_in),
    //     .S_out(S_out)
    // );
    KECCAK_f dut (
        .A_in(A_in),
        .A_out(A_out)
    );

    integer x, y;

    // Test stimulus
    initial begin
        // Apply stimulus
        //S_in = 'h1F00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000008000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        //S_in = 'h000000000000001f_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_8000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000;
        A_in[0][0] = 'h000000000000001f;
        A_in[1][0] = 'h0000000000000000;
        A_in[2][0] = 'h0000000000000000;
        A_in[3][0] = 'h0000000000000000;
        A_in[4][0] = 'h0000000000000000;
        A_in[0][1] = 'h0000000000000000;
        A_in[1][1] = 'h0000000000000000;
        A_in[2][1] = 'h0000000000000000;
        A_in[3][1] = 'h0000000000000000;
        A_in[4][1] = 'h0000000000000000;
        A_in[0][2] = 'h0000000000000000;
        A_in[1][2] = 'h0000000000000000;
        A_in[2][2] = 'h0000000000000000;
        A_in[3][2] = 'h0000000000000000;
        A_in[4][2] = 'h0000000000000000;
        A_in[0][3] = 'h0000000000000000;
        A_in[1][3] = 'h8000000000000000;
        A_in[2][3] = 'h0000000000000000;
        A_in[3][3] = 'h0000000000000000;
        A_in[4][3] = 'h0000000000000000;
        A_in[0][4] = 'h0000000000000000;
        A_in[1][4] = 'h0000000000000000;
        A_in[2][4] = 'h0000000000000000;
        A_in[3][4] = 'h0000000000000000;
        A_in[4][4] = 'h0000000000000000;
        
        // Wait for a few clock cycles
        #10;
        
        // Print the output
        // $display("S_in  =   %h", S_in);
        // $display("S_out =   %h", S_out);
        // $display("Expected: 1E000000000000001F00000000000000000000000000008000000000000000003E0000000000000001000000000000001F00000000000000000000000000008000000000000000003E0000000000000001000000000000001F00000000000000000000000000008000000000000000003E0000000000000001000000000000001F00000000000080000000000000008000000000000000003E0000000000000001000000000000001F00000000000000000000000000008000000000000000003E00000000000000");
        for (y = 0; y < 5; y = y + 1) begin
            for (x = 0; x < 5; x = x + 1) begin
                $display("A_in [%0d, %0d] = %h", x, y, A_in[x][y]);
            end
        end

        for (y = 0; y < 5; y = y + 1) begin
            for (x = 0; x < 5; x = x + 1) begin
                $display("A_out[%0d, %0d] = %h", x, y, A_out[x][y]);
            end
        end

        $display("Expected:");
        $display("A_out[0, 0] = 000000000000001e");
        $display("A_out[1, 0] = 000000000000001f");
        $display("A_out[2, 0] = 8000000000000000");
        $display("A_out[3, 0] = 0000000000000000");
        $display("A_out[4, 0] = 000000000000003e");
        $display("A_out[0, 1] = 0000000000000001");
        $display("A_out[1, 1] = 000000000000001f");
        $display("A_out[2, 1] = 8000000000000000");
        $display("A_out[3, 1] = 0000000000000000");
        $display("A_out[4, 1] = 000000000000003e");
        $display("A_out[0, 2] = 0000000000000001");
        $display("A_out[1, 2] = 000000000000001f");
        $display("A_out[2, 2] = 8000000000000000");
        $display("A_out[3, 2] = 0000000000000000");
        $display("A_out[4, 2] = 000000000000003e");
        $display("A_out[0, 3] = 0000000000000001");
        $display("A_out[1, 3] = 800000000000001f");
        $display("A_out[2, 3] = 8000000000000000");
        $display("A_out[3, 3] = 0000000000000000");
        $display("A_out[4, 3] = 000000000000003e");
        $display("A_out[0, 4] = 0000000000000001");
        $display("A_out[1, 4] = 000000000000001f");
        $display("A_out[2, 4] = 8000000000000000");
        $display("A_out[3, 4] = 0000000000000000");
        $display("A_out[4, 4] = 000000000000003e");

        // End the simulation
        $stop;
    end
    
endmodule
module SHAKE256_tb;



endmodule
`timescale 1ps/1ps

module KECCAK_f_tb;

    logic [1599:0] S_in, S_out;
    
    KECCAK_f dut (.S_in(S_in), .S_out(S_out));

    initial begin
        $dumpfile("KECCAKf_tb.vcd");
        $dumpvars;

        S_in = 'h1F00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000008000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        
        #1;
        
        $display("S_in  = %h", S_in);
        $display("S_out = %h", S_out);

        $finish;
    end
    
endmodule
module control_unit (
    input clock, reset,
    input [10:0] length,
    output [2:0] addrA, addrB,
    output [1:0] state_sel,
    output wren, busy, full, aclr, squeeze
);



endmodule